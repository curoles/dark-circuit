/* Core Debug Port (CDP).
 *
 * Authors: Igor Lesik 2021
 *
 * Core Debug Port makes the communation channel
 * between JTAG and Core Debug logic.
 *
 * CDP has two interfaces:
 *
 * - JTAG interface and
 * - memory bus interface to Core Debug logic..
 */
module CoreDbgPort (
);


endmodule: CoreDbgPort
