module TbTop (

);

    JtagTap _tap();

endmodule: TbTop
