module TbTop (

);

    localparam WIDTH = 64;

endmodule: TbTop
