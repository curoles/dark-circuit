module TbTop (

);

    DbgAccPort _dap();

endmodule: TbTop
