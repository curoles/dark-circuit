module TbTop (

);

endmodule: TbTop
