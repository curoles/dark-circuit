/*
 *
 *
 * http://bibl.ica.jku.at/dc/build/html/basiccircuits/basiccircuits.html
 *
 *
 */
